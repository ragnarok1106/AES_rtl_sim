module AES_TOP (
);

endmodule
