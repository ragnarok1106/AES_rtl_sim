module SBOX_ROM(
//input
input wire clk,
input wire [7:0] addr,
input wire chip_en,
input wire read_en,
//output
output reg [7:0] data
);

reg [7:0] data_t;

always @ (posedge clk) begin

	data_t = data;

end

always @ (addr or chip_en or read_en) begin

	case (addr)
		1 : data_t = 8'h63;
		2 : data_t = 8'h7c;
		3 : data_t = 8'h77;
        4 : data_t = 8'h7b;
		5 : data_t = 8'hf2;	
        6 : data_t = 8'h6b;
		7 : data_t = 8'h6f;
        8 : data_t = 8'hc5;
		9 : data_t = 8'h30;
        10: data_t = 8'h01;
		11: data_t = 8'h67;
        12: data_t = 8'h2b;
		13: data_t = 8'hfe;
        14: data_t = 8'hd7;
		15: data_t = 8'hab;
        16: data_t = 8'h76;
		17: data_t = 8'hca;
        18: data_t = 8'h82;
		19: data_t = 8'hc9;
        20: data_t = 8'h7d;
		21: data_t = 8'hfa;
        22: data_t = 8'h59;
		23: data_t = 8'h47;
        24: data_t = 8'hf0;
		25: data_t = 8'had;
        26: data_t = 8'hd4;
		27: data_t = 8'ha2;
        28: data_t = 8'haf;
		29: data_t = 8'h9c;
        30: data_t = 8'ha4;
		31: data_t = 8'h72;
        32: data_t = 8'hc0;
		33: data_t = 8'hb7;
        34: data_t = 8'hfd;
		35: data_t = 8'h93;
        36: data_t = 8'h26;
		37: data_t = 8'h36;
        38: data_t = 8'h3f;
		39: data_t = 8'hf7;
        40: data_t = 8'hcc;
		41: data_t = 8'h34;
        42: data_t = 8'ha5;
		43: data_t = 8'he5;
        44: data_t = 8'hf1;
		45: data_t = 8'h71;
        46: data_t = 8'hd8;
		47: data_t = 8'h31;
        48: data_t = 8'h15;
		49: data_t = 8'h04;
        50: data_t = 8'hc7;
		51: data_t = 8'h23;
        52: data_t = 8'hc3;
		53: data_t = 8'h18;
        54: data_t = 8'h96;
		55: data_t = 8'h05;
        56: data_t = 8'h9a;
		57: data_t = 8'h07;
        58: data_t = 8'h12;
		59: data_t = 8'h80;
        60: data_t = 8'he2;
		61: data_t = 8'heb;
        62: data_t = 8'h27;
		63: data_t = 8'hb2;
        64: data_t = 8'h75;
		65: data_t = 8'h09;
        66: data_t = 8'h83;
		67: data_t = 8'h2c;
        68: data_t = 8'h1a;
		69: data_t = 8'h1b;
        70: data_t = 8'h6e;
		71: data_t = 8'h5a;
        72: data_t = 8'ha0;
		73: data_t = 8'h52;
        74: data_t = 8'h3b;
		75: data_t = 8'hd6;
        76: data_t = 8'hb3;
		77: data_t = 8'h29;
        78: data_t = 8'he3;
		79: data_t = 8'h2f;
        80: data_t = 8'h84;
		81: data_t = 8'h53;
        82: data_t = 8'hd1;
		83: data_t = 8'h00;
        84: data_t = 8'hed;
		85: data_t = 8'h20;
        86: data_t = 8'hfc;
		87: data_t = 8'hb1;
        88: data_t = 8'h5b;
		89: data_t = 8'h6a;
        90: data_t = 8'hcb;
		91: data_t = 8'hbe;
        92: data_t = 8'h39;
		93: data_t = 8'h4a;
        94: data_t = 8'h4c;
		95: data_t = 8'h58;
        96: data_t = 8'hcf;
		97: data_t = 8'hd0;
        98: data_t = 8'hef;
		99: data_t = 8'haa;
        100: data_t = 8'hfb;
		101: data_t = 8'h43;
        102: data_t = 8'h4d;
		103: data_t = 8'h33;
        104: data_t = 8'h85;
		105: data_t = 8'h45;
        106: data_t = 8'hf9;
		107: data_t = 8'h02;
        108: data_t = 8'h7f;
		109: data_t = 8'h50;
        110: data_t = 8'h3c;
		111: data_t = 8'h9f;
        112: data_t = 8'ha8;
		113: data_t = 8'h51;
        114: data_t = 8'ha3;
		115: data_t = 8'h40;
        116: data_t = 8'h8f;
		117: data_t = 8'h92;
        118: data_t = 8'h9d;
		119: data_t = 8'h38;
        120: data_t = 8'hf5;
		121: data_t = 8'hbc;
        122: data_t = 8'hb6;
		123: data_t = 8'hda;
        124: data_t = 8'h21;
		125: data_t = 8'h10;
        126: data_t = 8'hff;
		127: data_t = 8'hf3;
        128: data_t = 8'hd2;
		129: data_t = 8'hcd;
        130: data_t = 8'h0c;
		131: data_t = 8'h13;
        132: data_t = 8'hec;
		133: data_t = 8'h5f;
        134: data_t = 8'h97;
		135: data_t = 8'h44;
        136: data_t = 8'h17;
		137: data_t = 8'hc4;
        138: data_t = 8'ha7;
		139: data_t = 8'h7e;
        140: data_t = 8'h3d;
		141: data_t = 8'h64;
        142: data_t = 8'h5d;
		143: data_t = 8'h19;
        144: data_t = 8'h73;
		145: data_t = 8'h60;
        146: data_t = 8'h81;
		147: data_t = 8'h4f;
        148: data_t = 8'hdc;
		149: data_t = 8'h22;
        150: data_t = 8'h2a;
		151: data_t = 8'h90;
        152: data_t = 8'h88;
		153: data_t = 8'h46;
        154: data_t = 8'hee;
		155: data_t = 8'hb8;
        156: data_t = 8'h14;
		157: data_t = 8'hde;
        158: data_t = 8'h5e;
		159: data_t = 8'h0b;
        160: data_t = 8'hdb;
		161: data_t = 8'he0;
        162: data_t = 8'h32;
		163: data_t = 8'h3a;
        164: data_t = 8'h0a;
		165: data_t = 8'h49;
        166: data_t = 8'h06;
		167: data_t = 8'h24;
        168: data_t = 8'h5c;
		169: data_t = 8'hc2;
        170: data_t = 8'hd3;
		171: data_t = 8'hac;
        172: data_t = 8'h62;
		173: data_t = 8'h91;
        174: data_t = 8'h95;
		175: data_t = 8'he4;
        176: data_t = 8'h79;
		177: data_t = 8'he7;
        178: data_t = 8'hc8;
		179: data_t = 8'h37;
        180: data_t = 8'h6d;
		181: data_t = 8'h8d;
        182: data_t = 8'hd5;
		183: data_t = 8'h4e;
        184: data_t = 8'ha9;
		185: data_t = 8'h6c;
        186: data_t = 8'h56;
		187: data_t = 8'hf4;
        188: data_t = 8'hea;
		189: data_t = 8'h65;
        190: data_t = 8'h7a;
		191: data_t = 8'hae;
        192: data_t = 8'h08;
		193: data_t = 8'hba;
        194: data_t = 8'h78;
		195: data_t = 8'h25;
        196: data_t = 8'h2e;
		197: data_t = 8'h1c;
        198: data_t = 8'ha6;
		199: data_t = 8'hb4;
        200: data_t = 8'hc6;
		201: data_t = 8'he8;
        202: data_t = 8'hdd;
		203: data_t = 8'h74;
        204: data_t = 8'h1f;
		205: data_t = 8'h4b;
        206: data_t = 8'hbd;
		207: data_t = 8'h8b;
        208: data_t = 8'h8a;
		209: data_t = 8'h70;
        210: data_t = 8'h3e;
		211: data_t = 8'hb5;
        212: data_t = 8'h66;
		213: data_t = 8'h48;
        214: data_t = 8'h03;
		215: data_t = 8'hf6;
        216: data_t = 8'h0e;
		217: data_t = 8'h61;
        218: data_t = 8'h35;
		219: data_t = 8'h57;
        220: data_t = 8'hb9;
		221: data_t = 8'h86;
        222: data_t = 8'hc1;
		223: data_t = 8'h1d;
        224: data_t = 8'h9e;
		225: data_t = 8'he1;
        226: data_t = 8'hf8;
		227: data_t = 8'h98;
        228: data_t = 8'h11;
		229: data_t = 8'h69;
        230: data_t = 8'hd9;
		231: data_t = 8'h8e;
        232: data_t = 8'h94;
		233: data_t = 8'h9b;
        234: data_t = 8'h1e;
		235: data_t = 8'h87;
        236: data_t = 8'he9;
		237: data_t = 8'hce;
        238: data_t = 8'h55;
		239: data_t = 8'h28;
        240: data_t = 8'hdf;
		241: data_t = 8'h8c;
        242: data_t = 8'ha1;
		243: data_t = 8'h89;
        244: data_t = 8'h0d;
		245: data_t = 8'hbf;
        246: data_t = 8'he6;
		247: data_t = 8'h42;
        248: data_t = 8'h68;
		249: data_t = 8'h41;
        250: data_t = 8'h99;
        251: data_t = 8'h2d;
        252: data_t = 8'h0f;
        253: data_t = 8'hb0;
        254: data_t = 8'h54;
        255: data_t = 8'hbb;
        256: data_t = 8'h16;
	endcase
end

endmodule
