module sbox_rom(
//input
input wire clk,
input wire [7:0] addr,
input wire chip_en,
input wire read_en,
//output
output reg [7:0] data
);

reg [7:0] data_t;

always @ (negedge clk) begin

	data = data_t;

end

always @ (addr or chip_en or read_en) begin

	case (addr)
		 0 : data_t = 8'h63;
		 1 : data_t = 8'h7c;
		 2 : data_t = 8'h77;
         3 : data_t = 8'h7b;
		 4 : data_t = 8'hf2;	
         5 : data_t = 8'h6b;
		 6 : data_t = 8'h6f;
         7 : data_t = 8'hc5;
		 8 : data_t = 8'h30;
         9 : data_t = 8'h01;
		 10: data_t = 8'h67;
         11: data_t = 8'h2b;
		 12: data_t = 8'hfe;
         13: data_t = 8'hd7;
		 14: data_t = 8'hab;
         15: data_t = 8'h76;
		 16: data_t = 8'hca;
         17: data_t = 8'h82;
		 18: data_t = 8'hc9;
         19: data_t = 8'h7d;
		 20: data_t = 8'hfa;
         21: data_t = 8'h59;
		 22: data_t = 8'h47;
         23: data_t = 8'hf0;
		 24: data_t = 8'had;
         25: data_t = 8'hd4;
		 26: data_t = 8'ha2;
         27: data_t = 8'haf;
		 28: data_t = 8'h9c;
         29: data_t = 8'ha4;
		 30: data_t = 8'h72;
         31: data_t = 8'hc0;
		 32: data_t = 8'hb7;
         33: data_t = 8'hfd;
		 34: data_t = 8'h93;
         35: data_t = 8'h26;
		 36: data_t = 8'h36;
         37: data_t = 8'h3f;
		 38: data_t = 8'hf7;
         39: data_t = 8'hcc;
		 40: data_t = 8'h34;
         41: data_t = 8'ha5;
		 42: data_t = 8'he5;
         43: data_t = 8'hf1;
		 44: data_t = 8'h71;
         45: data_t = 8'hd8;
		 46: data_t = 8'h31;
         47: data_t = 8'h15;
		 48: data_t = 8'h04;
         49: data_t = 8'hc7;
		 50: data_t = 8'h23;
         51: data_t = 8'hc3;
		 52: data_t = 8'h18;
         53: data_t = 8'h96;
		 54: data_t = 8'h05;
         55: data_t = 8'h9a;
		 56: data_t = 8'h07;
         57: data_t = 8'h12;
		 58: data_t = 8'h80;
         59: data_t = 8'he2;
		 60: data_t = 8'heb;
         61: data_t = 8'h27;
		 62: data_t = 8'hb2;
         63: data_t = 8'h75;
		 64: data_t = 8'h09;
         65: data_t = 8'h83;
		 66: data_t = 8'h2c;
         67: data_t = 8'h1a;
		 68: data_t = 8'h1b;
         69: data_t = 8'h6e;
		 70: data_t = 8'h5a;
         71: data_t = 8'ha0;
		 72: data_t = 8'h52;
         73: data_t = 8'h3b;
		 74: data_t = 8'hd6;
         75: data_t = 8'hb3;
		 76: data_t = 8'h29;
         77: data_t = 8'he3;
		 78: data_t = 8'h2f;
         79: data_t = 8'h84;
		 80: data_t = 8'h53;
         81: data_t = 8'hd1;
		 82: data_t = 8'h00;
         83: data_t = 8'hed;
		 84: data_t = 8'h20;
         85: data_t = 8'hfc;
		 86: data_t = 8'hb1;
         87: data_t = 8'h5b;
		 88: data_t = 8'h6a;
         89: data_t = 8'hcb;
		 90: data_t = 8'hbe;
         91: data_t = 8'h39;
		 92: data_t = 8'h4a;
         93: data_t = 8'h4c;
		 94: data_t = 8'h58;
         95: data_t = 8'hcf;
		 96: data_t = 8'hd0;
         97: data_t = 8'hef;
		 98: data_t = 8'haa;
         99: data_t = 8'hfb;
		 100: data_t = 8'h43;
         101: data_t = 8'h4d;
		 102: data_t = 8'h33;
         103: data_t = 8'h85;
		 104: data_t = 8'h45;
         105: data_t = 8'hf9;
		 106: data_t = 8'h02;
         107: data_t = 8'h7f;
		 108: data_t = 8'h50;
         109: data_t = 8'h3c;
		 110: data_t = 8'h9f;
         111: data_t = 8'ha8;
		 112: data_t = 8'h51;
         113: data_t = 8'ha3;
		 114: data_t = 8'h40;
         115: data_t = 8'h8f;
		 116: data_t = 8'h92;
         117: data_t = 8'h9d;
		 118: data_t = 8'h38;
         119: data_t = 8'hf5;
		 120: data_t = 8'hbc;
         121: data_t = 8'hb6;
		 122: data_t = 8'hda;
         123: data_t = 8'h21;
		 124: data_t = 8'h10;
         125: data_t = 8'hff;
		 126: data_t = 8'hf3;
         127: data_t = 8'hd2;
		 128: data_t = 8'hcd;
         129: data_t = 8'h0c;
		 130: data_t = 8'h13;
         131: data_t = 8'hec;
		 132: data_t = 8'h5f;
         133: data_t = 8'h97;
		 134: data_t = 8'h44;
         135: data_t = 8'h17;
		 136: data_t = 8'hc4;
         137: data_t = 8'ha7;
		 138: data_t = 8'h7e;
         139: data_t = 8'h3d;
		 140: data_t = 8'h64;
         141: data_t = 8'h5d;
		 142: data_t = 8'h19;
         143: data_t = 8'h73;
		 144: data_t = 8'h60;
         145: data_t = 8'h81;
		 146: data_t = 8'h4f;
         147: data_t = 8'hdc;
		 148: data_t = 8'h22;
         149: data_t = 8'h2a;
		 150: data_t = 8'h90;
         151: data_t = 8'h88;
		 152: data_t = 8'h46;
         153: data_t = 8'hee;
		 154: data_t = 8'hb8;
         155: data_t = 8'h14;
		 156: data_t = 8'hde;
         157: data_t = 8'h5e;
		 158: data_t = 8'h0b;
         159: data_t = 8'hdb;
		 160: data_t = 8'he0;
         161: data_t = 8'h32;
		 162: data_t = 8'h3a;
         163: data_t = 8'h0a;
		 164: data_t = 8'h49;
         165: data_t = 8'h06;
		 166: data_t = 8'h24;
         167: data_t = 8'h5c;
		 168: data_t = 8'hc2;
         169: data_t = 8'hd3;
		 170: data_t = 8'hac;
         171: data_t = 8'h62;
		 172: data_t = 8'h91;
         173: data_t = 8'h95;
		 174: data_t = 8'he4;
         175: data_t = 8'h79;
		 176: data_t = 8'he7;
         177: data_t = 8'hc8;
		 178: data_t = 8'h37;
         179: data_t = 8'h6d;
		 180: data_t = 8'h8d;
         181: data_t = 8'hd5;
		 182: data_t = 8'h4e;
         183: data_t = 8'ha9;
		 184: data_t = 8'h6c;
         185: data_t = 8'h56;
		 186: data_t = 8'hf4;
         187: data_t = 8'hea;
		 188: data_t = 8'h65;
         189: data_t = 8'h7a;
		 190: data_t = 8'hae;
         191: data_t = 8'h08;
		 192: data_t = 8'hba;
         193: data_t = 8'h78;
		 194: data_t = 8'h25;
         195: data_t = 8'h2e;
		 196: data_t = 8'h1c;
         197: data_t = 8'ha6;
		 198: data_t = 8'hb4;
         199: data_t = 8'hc6;
		 200: data_t = 8'he8;
         201: data_t = 8'hdd;
		 202: data_t = 8'h74;
         203: data_t = 8'h1f;
		 204: data_t = 8'h4b;
         205: data_t = 8'hbd;
		 206: data_t = 8'h8b;
         207: data_t = 8'h8a;
		 208: data_t = 8'h70;
         209: data_t = 8'h3e;
		 210: data_t = 8'hb5;
         211: data_t = 8'h66;
		 212: data_t = 8'h48;
         213: data_t = 8'h03;
		 214: data_t = 8'hf6;
         215: data_t = 8'h0e;
		 216: data_t = 8'h61;
         217: data_t = 8'h35;
		 218: data_t = 8'h57;
         219: data_t = 8'hb9;
		 220: data_t = 8'h86;
         221: data_t = 8'hc1;
		 222: data_t = 8'h1d;
         223: data_t = 8'h9e;
		 224: data_t = 8'he1;
         225: data_t = 8'hf8;
		 226: data_t = 8'h98;
         227: data_t = 8'h11;
		 228: data_t = 8'h69;
         229: data_t = 8'hd9;
		 230: data_t = 8'h8e;
         231: data_t = 8'h94;
		 232: data_t = 8'h9b;
         233: data_t = 8'h1e;
		 234: data_t = 8'h87;
         235: data_t = 8'he9;
		 236: data_t = 8'hce;
         237: data_t = 8'h55;
		 238: data_t = 8'h28;
         239: data_t = 8'hdf;
		 240: data_t = 8'h8c;
         241: data_t = 8'ha1;
		 242: data_t = 8'h89;
         243: data_t = 8'h0d;
		 244: data_t = 8'hbf;
         245: data_t = 8'he6;
		 246: data_t = 8'h42;
         247: data_t = 8'h68;
		 248: data_t = 8'h41;
         249: data_t = 8'h99;
         250: data_t = 8'h2d;
         251: data_t = 8'h0f;
         252: data_t = 8'hb0;
         253: data_t = 8'h54;
         254: data_t = 8'hbb;
         255: data_t = 8'h16;
	endcase
end

endmodule
